library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"417f7f00",
     1 => x"01000041",
     2 => x"180c0603",
     3 => x"00406030",
     4 => x"7f414100",
     5 => x"0800007f",
     6 => x"0603060c",
     7 => x"8000080c",
     8 => x"80808080",
     9 => x"00008080",
    10 => x"07030000",
    11 => x"00000004",
    12 => x"54547420",
    13 => x"0000787c",
    14 => x"44447f7f",
    15 => x"0000387c",
    16 => x"44447c38",
    17 => x"00000044",
    18 => x"44447c38",
    19 => x"00007f7f",
    20 => x"54547c38",
    21 => x"0000185c",
    22 => x"057f7e04",
    23 => x"00000005",
    24 => x"a4a4bc18",
    25 => x"00007cfc",
    26 => x"04047f7f",
    27 => x"0000787c",
    28 => x"7d3d0000",
    29 => x"00000040",
    30 => x"fd808080",
    31 => x"0000007d",
    32 => x"38107f7f",
    33 => x"0000446c",
    34 => x"7f3f0000",
    35 => x"7c000040",
    36 => x"0c180c7c",
    37 => x"0000787c",
    38 => x"04047c7c",
    39 => x"0000787c",
    40 => x"44447c38",
    41 => x"0000387c",
    42 => x"2424fcfc",
    43 => x"0000183c",
    44 => x"24243c18",
    45 => x"0000fcfc",
    46 => x"04047c7c",
    47 => x"0000080c",
    48 => x"54545c48",
    49 => x"00002074",
    50 => x"447f3f04",
    51 => x"00000044",
    52 => x"40407c3c",
    53 => x"00007c7c",
    54 => x"60603c1c",
    55 => x"3c001c3c",
    56 => x"6030607c",
    57 => x"44003c7c",
    58 => x"3810386c",
    59 => x"0000446c",
    60 => x"60e0bc1c",
    61 => x"00001c3c",
    62 => x"5c746444",
    63 => x"0000444c",
    64 => x"773e0808",
    65 => x"00004141",
    66 => x"7f7f0000",
    67 => x"00000000",
    68 => x"3e774141",
    69 => x"02000808",
    70 => x"02030101",
    71 => x"7f000102",
    72 => x"7f7f7f7f",
    73 => x"08007f7f",
    74 => x"3e1c1c08",
    75 => x"7f7f7f3e",
    76 => x"1c3e3e7f",
    77 => x"0008081c",
    78 => x"7c7c1810",
    79 => x"00001018",
    80 => x"7c7c3010",
    81 => x"10001030",
    82 => x"78606030",
    83 => x"4200061e",
    84 => x"3c183c66",
    85 => x"78004266",
    86 => x"c6c26a38",
    87 => x"6000386c",
    88 => x"00600000",
    89 => x"0e006000",
    90 => x"5d5c5b5e",
    91 => x"4c711e0e",
    92 => x"bfddf9c2",
    93 => x"c04bc04d",
    94 => x"02ab741e",
    95 => x"a6c487c7",
    96 => x"c578c048",
    97 => x"48a6c487",
    98 => x"66c478c1",
    99 => x"ee49731e",
   100 => x"86c887df",
   101 => x"ef49e0c0",
   102 => x"a5c487ee",
   103 => x"f0496a4a",
   104 => x"c6f187f0",
   105 => x"c185cb87",
   106 => x"abb7c883",
   107 => x"87c7ff04",
   108 => x"264d2626",
   109 => x"264b264c",
   110 => x"4a711e4f",
   111 => x"5ae1f9c2",
   112 => x"48e1f9c2",
   113 => x"fe4978c7",
   114 => x"4f2687dd",
   115 => x"711e731e",
   116 => x"aab7c04a",
   117 => x"c287d303",
   118 => x"05bfded9",
   119 => x"4bc187c4",
   120 => x"4bc087c2",
   121 => x"5be2d9c2",
   122 => x"d9c287c4",
   123 => x"d9c25ae2",
   124 => x"c14abfde",
   125 => x"a2c0c19a",
   126 => x"87e8ec49",
   127 => x"bfc6d9c2",
   128 => x"ded9c248",
   129 => x"08fcb0bf",
   130 => x"87e9fe78",
   131 => x"c44a711e",
   132 => x"49721e66",
   133 => x"2687f3ea",
   134 => x"ff1e4f26",
   135 => x"ffc348d4",
   136 => x"48d0ff78",
   137 => x"ff78e1c0",
   138 => x"78c148d4",
   139 => x"30c44871",
   140 => x"7808d4ff",
   141 => x"c048d0ff",
   142 => x"4f2678e0",
   143 => x"5c5b5e0e",
   144 => x"86f40e5d",
   145 => x"c048a6c4",
   146 => x"bfec4b78",
   147 => x"ddf9c27e",
   148 => x"bfe84dbf",
   149 => x"ded9c24c",
   150 => x"f1e349bf",
   151 => x"49f7c187",
   152 => x"7087f5e6",
   153 => x"87d50298",
   154 => x"bfded9c2",
   155 => x"87dee349",
   156 => x"f7c14bc1",
   157 => x"87e0e649",
   158 => x"eb059870",
   159 => x"029b7387",
   160 => x"c287fac0",
   161 => x"05bfc6d9",
   162 => x"a6c887c7",
   163 => x"c578c148",
   164 => x"48a6c887",
   165 => x"d9c278c0",
   166 => x"66c848c6",
   167 => x"1efcca78",
   168 => x"c90266cc",
   169 => x"48a6cc87",
   170 => x"78d9d7c2",
   171 => x"a6cc87c7",
   172 => x"e4d7c248",
   173 => x"4966cc78",
   174 => x"c487f5cc",
   175 => x"cb4bc086",
   176 => x"e1ce49ee",
   177 => x"58a6cc87",
   178 => x"cbe549c7",
   179 => x"05987087",
   180 => x"496e87c8",
   181 => x"c10299c1",
   182 => x"4bc187c3",
   183 => x"c27ebfec",
   184 => x"49bfded9",
   185 => x"c887e7e1",
   186 => x"c5ce4966",
   187 => x"02987087",
   188 => x"d9c287d8",
   189 => x"c149bfc2",
   190 => x"c6d9c2b9",
   191 => x"d9fc7159",
   192 => x"49eecb87",
   193 => x"cc87dfcd",
   194 => x"49c758a6",
   195 => x"7087c9e4",
   196 => x"c5ff0598",
   197 => x"c1496e87",
   198 => x"fdfe0599",
   199 => x"029b7387",
   200 => x"49ff87d0",
   201 => x"c187e5fa",
   202 => x"ebe349da",
   203 => x"48a6c487",
   204 => x"d9c278c1",
   205 => x"c105bfde",
   206 => x"d9c287e2",
   207 => x"c002bfc6",
   208 => x"a6c487f1",
   209 => x"c0c0c848",
   210 => x"cad9c278",
   211 => x"bf976e7e",
   212 => x"c1486e49",
   213 => x"717e7080",
   214 => x"7087fde2",
   215 => x"c3c00298",
   216 => x"b466c487",
   217 => x"c14866c4",
   218 => x"a6c828b7",
   219 => x"05987058",
   220 => x"c387daff",
   221 => x"dfe249fd",
   222 => x"49fac387",
   223 => x"7487d9e2",
   224 => x"99ffc349",
   225 => x"49c01e71",
   226 => x"7487c1fa",
   227 => x"29b7c849",
   228 => x"49c11e71",
   229 => x"c887f5f9",
   230 => x"87f8c886",
   231 => x"ffc34974",
   232 => x"2cb7c899",
   233 => x"9c74b471",
   234 => x"87e0c002",
   235 => x"bfdad9c2",
   236 => x"87feca49",
   237 => x"c0059870",
   238 => x"4cc087c5",
   239 => x"c287d3c0",
   240 => x"e1ca49e0",
   241 => x"ded9c287",
   242 => x"87c6c058",
   243 => x"48dad9c2",
   244 => x"497478c0",
   245 => x"c00599c2",
   246 => x"ebc387ce",
   247 => x"87f8e049",
   248 => x"99c24970",
   249 => x"87cec002",
   250 => x"4aa5d8c1",
   251 => x"c5c0026a",
   252 => x"49fb4b87",
   253 => x"49740f73",
   254 => x"c00599c1",
   255 => x"f4c387ce",
   256 => x"87d4e049",
   257 => x"99c24970",
   258 => x"87cfc002",
   259 => x"7ea5d8c1",
   260 => x"c002bf6e",
   261 => x"fa4b87c5",
   262 => x"740f7349",
   263 => x"0599c849",
   264 => x"c387cfc0",
   265 => x"dfff49f5",
   266 => x"497087ee",
   267 => x"c00299c2",
   268 => x"f9c287e6",
   269 => x"c002bfe1",
   270 => x"c14887ca",
   271 => x"e5f9c288",
   272 => x"87cfc058",
   273 => x"7ea5d8c1",
   274 => x"c002bf6e",
   275 => x"ff4b87c5",
   276 => x"c40f7349",
   277 => x"78c148a6",
   278 => x"99c44974",
   279 => x"87cfc005",
   280 => x"ff49f2c3",
   281 => x"7087f1de",
   282 => x"0299c249",
   283 => x"c287ecc0",
   284 => x"7ebfe1f9",
   285 => x"a8b7c748",
   286 => x"87cbc003",
   287 => x"80c1486e",
   288 => x"58e5f9c2",
   289 => x"c187cfc0",
   290 => x"6e7ea5d8",
   291 => x"c5c002bf",
   292 => x"49fe4b87",
   293 => x"a6c40f73",
   294 => x"c378c148",
   295 => x"ddff49fd",
   296 => x"497087f6",
   297 => x"c00299c2",
   298 => x"f9c287e5",
   299 => x"c002bfe1",
   300 => x"f9c287c9",
   301 => x"78c048e1",
   302 => x"c187cfc0",
   303 => x"6e7ea5d8",
   304 => x"c5c002bf",
   305 => x"49fd4b87",
   306 => x"a6c40f73",
   307 => x"c378c148",
   308 => x"ddff49fa",
   309 => x"497087c2",
   310 => x"c00299c2",
   311 => x"f9c287e9",
   312 => x"c748bfe1",
   313 => x"c003a8b7",
   314 => x"f9c287c9",
   315 => x"78c748e1",
   316 => x"c187cfc0",
   317 => x"6e7ea5d8",
   318 => x"c5c002bf",
   319 => x"49fc4b87",
   320 => x"a6c40f73",
   321 => x"c078c148",
   322 => x"dcf9c24b",
   323 => x"cb50c048",
   324 => x"d1c549ee",
   325 => x"58a6cc87",
   326 => x"97dcf9c2",
   327 => x"dec105bf",
   328 => x"c3497487",
   329 => x"c00599f0",
   330 => x"dac187cd",
   331 => x"e7dbff49",
   332 => x"02987087",
   333 => x"c187c8c1",
   334 => x"4cbfe84b",
   335 => x"99ffc349",
   336 => x"712cb7c8",
   337 => x"ded9c2b4",
   338 => x"d8ff49bf",
   339 => x"66c887c0",
   340 => x"87dec449",
   341 => x"c0029870",
   342 => x"f9c287c6",
   343 => x"50c148dc",
   344 => x"97dcf9c2",
   345 => x"d6c005bf",
   346 => x"c3497487",
   347 => x"ff0599f0",
   348 => x"dac187c5",
   349 => x"dfdaff49",
   350 => x"05987087",
   351 => x"7387f8fe",
   352 => x"dcc0029b",
   353 => x"48a6c887",
   354 => x"bfe1f9c2",
   355 => x"4966c878",
   356 => x"a17591cb",
   357 => x"02bf6e7e",
   358 => x"4b87c6c0",
   359 => x"734966c8",
   360 => x"0266c40f",
   361 => x"c287c8c0",
   362 => x"49bfe1f9",
   363 => x"c287f8ee",
   364 => x"02bfe2d9",
   365 => x"4987ddc0",
   366 => x"7087f7c2",
   367 => x"d3c00298",
   368 => x"e1f9c287",
   369 => x"deee49bf",
   370 => x"ef49c087",
   371 => x"d9c287fe",
   372 => x"78c048e2",
   373 => x"d8ef8ef4",
   374 => x"796f4a87",
   375 => x"7379656b",
   376 => x"006e6f20",
   377 => x"6b796f4a",
   378 => x"20737965",
   379 => x"0066666f",
   380 => x"5c5b5e0e",
   381 => x"711e0e5d",
   382 => x"ddf9c24c",
   383 => x"cdc149bf",
   384 => x"d1c14da1",
   385 => x"747e6981",
   386 => x"87cf029c",
   387 => x"744ba5c4",
   388 => x"ddf9c27b",
   389 => x"e0ee49bf",
   390 => x"747b6e87",
   391 => x"87c4059c",
   392 => x"87c24bc0",
   393 => x"49734bc1",
   394 => x"d487e1ee",
   395 => x"87c80266",
   396 => x"87f2c049",
   397 => x"87c24a70",
   398 => x"d9c24ac0",
   399 => x"ed265ae6",
   400 => x"000087ef",
   401 => x"00000000",
   402 => x"12580000",
   403 => x"1b1d1411",
   404 => x"595a231c",
   405 => x"f2f59491",
   406 => x"0000f4eb",
   407 => x"00000000",
   408 => x"00000000",
   409 => x"711e0000",
   410 => x"bfc8ff4a",
   411 => x"48a17249",
   412 => x"ff1e4f26",
   413 => x"fe89bfc8",
   414 => x"c0c0c0c0",
   415 => x"c401a9c0",
   416 => x"c24ac087",
   417 => x"724ac187",
   418 => x"0e4f2648",
   419 => x"5d5c5b5e",
   420 => x"ff4b710e",
   421 => x"66d04cd4",
   422 => x"d678c048",
   423 => x"efd7ff49",
   424 => x"7cffc387",
   425 => x"ffc3496c",
   426 => x"494d7199",
   427 => x"c199f0c3",
   428 => x"cb05a9e0",
   429 => x"7cffc387",
   430 => x"98c3486c",
   431 => x"780866d0",
   432 => x"6c7cffc3",
   433 => x"31c8494a",
   434 => x"6c7cffc3",
   435 => x"72b2714a",
   436 => x"c331c849",
   437 => x"4a6c7cff",
   438 => x"4972b271",
   439 => x"ffc331c8",
   440 => x"714a6c7c",
   441 => x"48d0ffb2",
   442 => x"7378e0c0",
   443 => x"87c2029b",
   444 => x"48757b72",
   445 => x"4c264d26",
   446 => x"4f264b26",
   447 => x"0e4f261e",
   448 => x"0e5c5b5e",
   449 => x"1e7686f8",
   450 => x"fd49a6c8",
   451 => x"86c487fd",
   452 => x"486e4b70",
   453 => x"c203a8c2",
   454 => x"4a7387f0",
   455 => x"c19af0c3",
   456 => x"c702aad0",
   457 => x"aae0c187",
   458 => x"87dec205",
   459 => x"99c84973",
   460 => x"ff87c302",
   461 => x"4c7387c6",
   462 => x"acc29cc3",
   463 => x"87c2c105",
   464 => x"c94966c4",
   465 => x"c41e7131",
   466 => x"92d44a66",
   467 => x"49e5f9c2",
   468 => x"c9fe8172",
   469 => x"49d887f1",
   470 => x"87f4d4ff",
   471 => x"c21ec0c8",
   472 => x"fd49cee8",
   473 => x"ff87f7e5",
   474 => x"e0c048d0",
   475 => x"cee8c278",
   476 => x"4a66cc1e",
   477 => x"f9c292d4",
   478 => x"817249e5",
   479 => x"87f9c7fe",
   480 => x"acc186cc",
   481 => x"87c2c105",
   482 => x"c94966c4",
   483 => x"c41e7131",
   484 => x"92d44a66",
   485 => x"49e5f9c2",
   486 => x"c8fe8172",
   487 => x"e8c287e9",
   488 => x"66c81ece",
   489 => x"c292d44a",
   490 => x"7249e5f9",
   491 => x"fac5fe81",
   492 => x"ff49d787",
   493 => x"c887d9d3",
   494 => x"e8c21ec0",
   495 => x"e3fd49ce",
   496 => x"86cc87f5",
   497 => x"c048d0ff",
   498 => x"8ef878e0",
   499 => x"0e87e7fc",
   500 => x"5d5c5b5e",
   501 => x"ff4a710e",
   502 => x"66d04cd4",
   503 => x"adb7c34d",
   504 => x"c087c506",
   505 => x"87e1c148",
   506 => x"4b751e72",
   507 => x"f9c293d4",
   508 => x"497383e5",
   509 => x"87c1c0fe",
   510 => x"4b6b83c8",
   511 => x"c848d0ff",
   512 => x"7cdd78e1",
   513 => x"ffc34873",
   514 => x"737c7098",
   515 => x"29b7c849",
   516 => x"ffc34871",
   517 => x"737c7098",
   518 => x"29b7d049",
   519 => x"ffc34871",
   520 => x"737c7098",
   521 => x"28b7d848",
   522 => x"7cc07c70",
   523 => x"7c7c7c7c",
   524 => x"7c7c7c7c",
   525 => x"ff7c7c7c",
   526 => x"e0c048d0",
   527 => x"dc1e7578",
   528 => x"f0d1ff49",
   529 => x"7386c887",
   530 => x"87e8fa48",
   531 => x"c44a711e",
   532 => x"f9c249a2",
   533 => x"786a48c8",
   534 => x"48c2d9c2",
   535 => x"d9c27869",
   536 => x"e649bfc2",
   537 => x"d1ff87f4",
   538 => x"4f2687fd",
   539 => x"c44a711e",
   540 => x"f9c249a2",
   541 => x"c27abfc8",
   542 => x"79bfc2d9",
   543 => x"711e4f26",
   544 => x"c0029a4a",
   545 => x"c21e87ee",
   546 => x"fd49c4f5",
   547 => x"c487eafd",
   548 => x"02987086",
   549 => x"e8c287de",
   550 => x"f5c21ece",
   551 => x"c2fe49c4",
   552 => x"86c487c9",
   553 => x"cb029870",
   554 => x"cee8c287",
   555 => x"87dcfe49",
   556 => x"87c248c1",
   557 => x"4f2648c0",
   558 => x"9a4a711e",
   559 => x"87eec002",
   560 => x"c4f5c21e",
   561 => x"f0fcfd49",
   562 => x"7086c487",
   563 => x"87de0298",
   564 => x"49cee8c2",
   565 => x"c287d5fe",
   566 => x"c21ecee8",
   567 => x"fe49c4f5",
   568 => x"c487d6c2",
   569 => x"02987086",
   570 => x"48c187c4",
   571 => x"48c087c2",
   572 => x"c11e4f26",
   573 => x"c048cce7",
   574 => x"cdfac250",
   575 => x"87cc05bf",
   576 => x"49ffe4c2",
   577 => x"87e1d5fe",
   578 => x"58d1fac2",
   579 => x"48cce7c1",
   580 => x"fac250c2",
   581 => x"cc05bfd1",
   582 => x"cbe5c287",
   583 => x"c8d5fe49",
   584 => x"d5fac287",
   585 => x"d5fac258",
   586 => x"87d105bf",
   587 => x"c21ef1c0",
   588 => x"fe49d7e5",
   589 => x"c487c5db",
   590 => x"d9fac286",
   591 => x"564f2658",
   592 => x"30324349",
   593 => x"52202020",
   594 => x"4d004d4f",
   595 => x"43414745",
   596 => x"52545241",
   597 => x"4d004d4f",
   598 => x"43414745",
   599 => x"4e545241",
   600 => x"1e002056",
   601 => x"4bc01e73",
   602 => x"48cdfac2",
   603 => x"fac278c0",
   604 => x"78c048d1",
   605 => x"48d5fac2",
   606 => x"f5fd78c0",
   607 => x"d1e7c287",
   608 => x"c4f5c21e",
   609 => x"f0f9fd49",
   610 => x"7086c487",
   611 => x"87c90298",
   612 => x"bfc8f5c2",
   613 => x"d0c2fe49",
   614 => x"87d6fd87",
   615 => x"c2fe49c0",
   616 => x"fac287c7",
   617 => x"cd02bfd1",
   618 => x"c8f9c287",
   619 => x"c0c848bf",
   620 => x"f9c2b0c0",
   621 => x"ccff58cc",
   622 => x"fac287ed",
   623 => x"c405bfcd",
   624 => x"dde7c287",
   625 => x"c448734b",
   626 => x"264d2687",
   627 => x"264b264c",
   628 => x"4148434f",
   629 => x"2030324d",
   630 => x"20202020",
   631 => x"4d4f5200",
   632 => x"69616620",
   633 => x"0064656c",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
